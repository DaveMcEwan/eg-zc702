
module pl_m (
  // clkrst
  input  wire       i_clk0,
  input  wire       i_clk1,
  input  wire       i_clk2,
  input  wire       i_clk3,
  input  wire       i_rst,
  input  wire       i_ic_rst,

  // {{{ AXI ports from PS7
  input  wire          i_M_AXI_GP0_ARVALID,
  input  wire          i_M_AXI_GP0_AWVALID,
  input  wire          i_M_AXI_GP0_BREADY,
  input  wire          i_M_AXI_GP0_RREADY,
  input  wire          i_M_AXI_GP0_WLAST,
  input  wire          i_M_AXI_GP0_WVALID,
  input  wire [11:0]   i_M_AXI_GP0_ARID,
  input  wire [11:0]   i_M_AXI_GP0_AWID,
  input  wire [11:0]   i_M_AXI_GP0_WID,
  input  wire [1:0]    i_M_AXI_GP0_ARBURST,
  input  wire [1:0]    i_M_AXI_GP0_ARLOCK,
  input  wire [2:0]    i_M_AXI_GP0_ARSIZE,
  input  wire [1:0]    i_M_AXI_GP0_AWBURST,
  input  wire [1:0]    i_M_AXI_GP0_AWLOCK,
  input  wire [2:0]    i_M_AXI_GP0_AWSIZE,
  input  wire [2:0]    i_M_AXI_GP0_ARPROT,
  input  wire [2:0]    i_M_AXI_GP0_AWPROT,
  input  wire [31:0]   i_M_AXI_GP0_ARADDR,
  input  wire [31:0]   i_M_AXI_GP0_AWADDR,
  input  wire [31:0]   i_M_AXI_GP0_WDATA,
  input  wire [3:0]    i_M_AXI_GP0_ARCACHE,
  input  wire [3:0]    i_M_AXI_GP0_ARLEN,
  input  wire [3:0]    i_M_AXI_GP0_ARQOS,
  input  wire [3:0]    i_M_AXI_GP0_AWCACHE,
  input  wire [3:0]    i_M_AXI_GP0_AWLEN,
  input  wire [3:0]    i_M_AXI_GP0_AWQOS,
  input  wire [3:0]    i_M_AXI_GP0_WSTRB,
  output wire          o_M_AXI_GP0_ARREADY,
  output wire          o_M_AXI_GP0_AWREADY,
  output wire          o_M_AXI_GP0_BVALID,
  output wire          o_M_AXI_GP0_RLAST,
  output wire          o_M_AXI_GP0_RVALID,
  output wire          o_M_AXI_GP0_WREADY,
  output wire [11:0]   o_M_AXI_GP0_BID,
  output wire [11:0]   o_M_AXI_GP0_RID,
  output wire [1:0]    o_M_AXI_GP0_BRESP,
  output wire [1:0]    o_M_AXI_GP0_RRESP,
  output wire [31:0]   o_M_AXI_GP0_RDATA,

  input  wire          i_M_AXI_GP1_ARVALID,
  input  wire          i_M_AXI_GP1_AWVALID,
  input  wire          i_M_AXI_GP1_BREADY,
  input  wire          i_M_AXI_GP1_RREADY,
  input  wire          i_M_AXI_GP1_WLAST,
  input  wire          i_M_AXI_GP1_WVALID,
  input  wire [11:0]   i_M_AXI_GP1_ARID,
  input  wire [11:0]   i_M_AXI_GP1_AWID,
  input  wire [11:0]   i_M_AXI_GP1_WID,
  input  wire [1:0]    i_M_AXI_GP1_ARBURST,
  input  wire [1:0]    i_M_AXI_GP1_ARLOCK,
  input  wire [2:0]    i_M_AXI_GP1_ARSIZE,
  input  wire [1:0]    i_M_AXI_GP1_AWBURST,
  input  wire [1:0]    i_M_AXI_GP1_AWLOCK,
  input  wire [2:0]    i_M_AXI_GP1_AWSIZE,
  input  wire [2:0]    i_M_AXI_GP1_ARPROT,
  input  wire [2:0]    i_M_AXI_GP1_AWPROT,
  input  wire [31:0]   i_M_AXI_GP1_ARADDR,
  input  wire [31:0]   i_M_AXI_GP1_AWADDR,
  input  wire [31:0]   i_M_AXI_GP1_WDATA,
  input  wire [3:0]    i_M_AXI_GP1_ARCACHE,
  input  wire [3:0]    i_M_AXI_GP1_ARLEN,
  input  wire [3:0]    i_M_AXI_GP1_ARQOS,
  input  wire [3:0]    i_M_AXI_GP1_AWCACHE,
  input  wire [3:0]    i_M_AXI_GP1_AWLEN,
  input  wire [3:0]    i_M_AXI_GP1_AWQOS,
  input  wire [3:0]    i_M_AXI_GP1_WSTRB,
  output wire          o_M_AXI_GP1_ARREADY,
  output wire          o_M_AXI_GP1_AWREADY,
  output wire          o_M_AXI_GP1_BVALID,
  output wire          o_M_AXI_GP1_RLAST,
  output wire          o_M_AXI_GP1_RVALID,
  output wire          o_M_AXI_GP1_WREADY,
  output wire [11:0]   o_M_AXI_GP1_BID,
  output wire [11:0]   o_M_AXI_GP1_RID,
  output wire [1:0]    o_M_AXI_GP1_BRESP,
  output wire [1:0]    o_M_AXI_GP1_RRESP,
  output wire [31:0]   o_M_AXI_GP1_RDATA,
  // }}}

  output wire [7:0] o_led
);

  assign o_led = 8'h55;

endmodule

